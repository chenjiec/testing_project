library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_textio.all;
use ieee.numeric_std.all;
use work.myTypes.all;
use work.all;

entity tb_dlx is
end tb_dlx;

architecture tb of tb_dlx is
component DLX is 
port(clk:in std_logic; 
     rst:in std_logic);
end component;
signal clk:std_logic;
signal rst:std_logic;
begin
p1:DLX
port map(clk,rst);
process
begin
rst<='1','0'after 5 ns;
wait for 5 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';wait for 1 ns;
clk<='0';
wait for 1 ns;
clk<='1';
wait;
end process;
end tb;