library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use work.myTypes.all;

entity RF_file is
port(clk:in std_logic;
     reg_num:in std_logic_vector(4 downto 0);
     mux_stage5_out:in std_logic_vector(31 downto 0);
     RF_WE  :in std_logic;
     IR_LATCH_EN:in std_logic;
     reg_val:out std_logic_vector(31 downto 0)
   );
end RF_file;

architecture behavior of RF_file is
type re_mem is array (integer range 0 to 31) of std_logic_vector(31 downto 0);
signal reg: re_mem :=( "00000000000000000000000000000000",
                       "00000000000000000000000000000001",
                       "00000000000000000000000000000010",
                       "00000000000000000000000000000011",
                        
                       "00000000000000000000000000000100",                         
                       "00000000000000000000000000000001",
                       "00000000000000000000000000000010",
                       "00000000000000000000000000000011",
                        
                       "00000000000000000000000000000100",
                       "00000000000000000000000000000001",
                       "00000000000000000000000000000010",
                       "00000000000000000000000000000011", 
                       
                       "00000000000000000000000000000100",                         
                       "00000000000000000000000000000001",
                       "00000000000000000000000000000010",
                       "00000000000000000000000000000011",
                        
                       "00000000000000000000000000000100",
                       "00000000000000000000000000000001",
                       "00000000000000000000000000000010",
                       "00000000000000000000000000000011",  
                       
                       "00000000000000000000000000000100",                         
                       "00000000000000000000000000000001",
                       "00000000000000000000000000000010",
                       "00000000000000000000000000000011",
                        
                       "00000000000000000000000000000100",
                       "00000000000000000000000000000001",
                       "00000000000000000000000000000010",
                       "00000000000000000000000000000011", 
                       
                       "00000000000000000000000000000100",                         
                       "00000000000000000000000000000001",
                       "00000000000000000000000000000010",
                       "00000000000000000000000000000011"
                     );
begin
process(RF_WE,IR_LATCH_EN,clk)
begin
if(clk='1' and clk'event) then
if(RF_WE='0')then
reg_val<=reg(conv_integer(reg_num));
else
reg(conv_integer(reg_num))<=mux_stage5_out;
end if;
end if;
end process;
end behavior;
                       